--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   18:14:23 02/19/2018
-- Design Name:   
-- Module Name:   C:/Users/Jet/Documents/GitHub/AdvancedLogicCircuitProject/advalog_project/trafficLightTB.vhd
-- Project Name:  advalog_project
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: Entity_TrafficLight
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY trafficLightTB IS
END trafficLightTB;
 
ARCHITECTURE behavior OF trafficLightTB IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT Entity_TrafficLight
    PORT(
         clk : IN  std_logic;
         clr : IN  std_logic;
         light : OUT  std_logic_vector(10 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal clk : std_logic := '0';
   signal clr : std_logic := '0';

 	--Outputs
   signal light : std_logic_vector(10 downto 0);

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: Entity_TrafficLight PORT MAP (
          clk => clk,
          clr => clr,
          light => light
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
	



      -- insert stimulus here 

      wait;
   end process;

END;
